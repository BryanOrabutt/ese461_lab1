
module problem5(rst, req_0, req_1, gnt_0, gnt_1, idle);

input rst, req_0, req_1;
output reg gnt_0, gnt_1, idle;



endmodule
